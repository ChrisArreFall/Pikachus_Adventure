module pokecoin(input logic [9:0] x,y,pos_x,pos_y,
				 input logic en,enable,
				 output logic [7:0] r,g,b);

				logic [1:0] pokecoin_static [0:31][0:31]  = 	'{
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
																			'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}
																			};


				always_comb
					if(enable)
						case(pokecoin_static[y-pos_y][x-pos_x-1])
							3'b000 : {b,g,r} = 24'hebce87;//0x00000000
							3'b001 : {b,g,r} = 24'h0decf4;//0xff0decf4
							3'b010 : {b,g,r} = 24'h000000;//0xff000000
							3'b011 : {b,g,r} = 24'h0000ff;//0xff0000ff
							3'b100 : {b,g,r} = 24'hDCF5F5;//0xffffffff
							default: {b,g,r} = 24'hebce87;
						endcase
					else
						{b,g,r} = 24'hebce87;

endmodule
