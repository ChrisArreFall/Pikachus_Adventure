module coin();




endmodule


