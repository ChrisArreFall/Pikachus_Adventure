module cloud();



endmodule
